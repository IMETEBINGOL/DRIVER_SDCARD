localparam      SPI_SPI_INTERFACE_PACKAGE_WIDTH     = 8;